module rom(addr,data);
	input [6:0] addr;
	output reg [15:0] data;
	
	//Look-up Table of Sigmoid (X >=0)
	always @ (addr) begin
		case(addr)
			7'b0 : data = 16'b10000000;
			7'b1 : data = 16'b10000100;
			7'b10 : data = 16'b10001000;
			7'b11 : data = 16'b10001100;
			7'b100 : data = 16'b10010000;
			7'b101 : data = 16'b10010100;
			7'b110 : data = 16'b10011000;
			7'b111 : data = 16'b10011100;
			7'b1000 : data = 16'b10011111;
			7'b1001 : data = 16'b10100011;
			7'b1010 : data = 16'b10100111;
			7'b1011 : data = 16'b10101010;
			7'b1100 : data = 16'b10101110;
			7'b1101 : data = 16'b10110001;
			7'b1110 : data = 16'b10110101;
			7'b1111 : data = 16'b10111000;
			7'b10000 : data = 16'b10111011;
			7'b10001 : data = 16'b10111110;
			7'b10010 : data = 16'b11000001;
			7'b10011 : data = 16'b11000100;
			7'b10100 : data = 16'b11000111;
			7'b10101 : data = 16'b11001010;
			7'b10110 : data = 16'b11001100;
			7'b10111 : data = 16'b11001111;
			7'b11000 : data = 16'b11010001;
			7'b11001 : data = 16'b11010100;
			7'b11010 : data = 16'b11010110;
			7'b11011 : data = 16'b11011000;
			7'b11100 : data = 16'b11011010;
			7'b11101 : data = 16'b11011100;
			7'b11110 : data = 16'b11011110;
			7'b11111 : data = 16'b11100000;
			7'b100000 : data = 16'b11100001;
			7'b100001 : data = 16'b11100011;
			7'b100010 : data = 16'b11100101;
			7'b100011 : data = 16'b11100110;
			7'b100100 : data = 16'b11101000;
			7'b100101 : data = 16'b11101001;
			7'b100110 : data = 16'b11101010;
			7'b100111 : data = 16'b11101011;
			7'b101000 : data = 16'b11101101;
			7'b101001 : data = 16'b11101110;
			7'b101010 : data = 16'b11101111;
			7'b101011 : data = 16'b11110000;
			7'b101100 : data = 16'b11110001;
			7'b101101 : data = 16'b11110001;
			7'b101110 : data = 16'b11110010;
			7'b101111 : data = 16'b11110011;
			7'b110000 : data = 16'b11110100;
			7'b110001 : data = 16'b11110101;
			7'b110010 : data = 16'b11110101;
			7'b110011 : data = 16'b11110110;
			7'b110100 : data = 16'b11110110;
			7'b110101 : data = 16'b11110111;
			7'b110110 : data = 16'b11111000;
			7'b110111 : data = 16'b11111000;
			7'b111000 : data = 16'b11111000;
			7'b111001 : data = 16'b11111001;
			7'b111010 : data = 16'b11111001;
			7'b111011 : data = 16'b11111010;
			7'b111100 : data = 16'b11111010;
			7'b111101 : data = 16'b11111010;
			7'b111110 : data = 16'b11111011;
			7'b111111 : data = 16'b11111011;
			7'b1000000 : data = 16'b11111011;
			7'b1000001 : data = 16'b11111100;
			7'b1000010 : data = 16'b11111100;
			7'b1000011 : data = 16'b11111100;
			7'b1000100 : data = 16'b11111100;
			7'b1000101 : data = 16'b11111101;
			7'b1000110 : data = 16'b11111101;
			7'b1000111 : data = 16'b11111101;
			7'b1001000 : data = 16'b11111101;
			7'b1001001 : data = 16'b11111101;
			7'b1001010 : data = 16'b11111110;
			7'b1001011 : data = 16'b11111110;
			7'b1001100 : data = 16'b11111110;
			7'b1001101 : data = 16'b11111110;
			7'b1001110 : data = 16'b11111110;
			7'b1001111 : data = 16'b11111110;
			7'b1010000 : data = 16'b11111110;
			7'b1010001 : data = 16'b11111110;
			7'b1010010 : data = 16'b11111110;
			7'b1010011 : data = 16'b11111111;
			7'b1010100 : data = 16'b11111111;
			7'b1010101 : data = 16'b11111111;
			7'b1010110 : data = 16'b11111111;
			7'b1010111 : data = 16'b11111111;
			7'b1011000 : data = 16'b11111111;
			7'b1011001 : data = 16'b11111111;
			7'b1011010 : data = 16'b11111111;
			7'b1011011 : data = 16'b11111111;
			7'b1011100 : data = 16'b11111111;
			7'b1011101 : data = 16'b11111111;
			7'b1011110 : data = 16'b11111111;
			7'b1011111 : data = 16'b11111111;
			7'b1100000 : data = 16'b11111111;
		endcase	
	end
	
endmodule
