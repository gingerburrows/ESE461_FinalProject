`timescale 1ns / 1ps
module rom(addr,data);
	input [15:0] addr;
	output reg [15:0] data;
	
	//Look-up Table of Sigmoid (X >=0)
	always @ (addr) begin
		case(addr)
			16'b0 : data = 16'b10000000;
			16'b11010 : data = 16'b10000110;
			16'b110011 : data = 16'b10001101;
			16'b1001101 : data = 16'b10010011;
			16'b1100110 : data = 16'b10011001;
			16'b10000000 : data = 16'b10011111;
			16'b10011010 : data = 16'b10100101;
			16'b10110011 : data = 16'b10101011;
			16'b11001101 : data = 16'b10110001;
			16'b11100110 : data = 16'b10110110;
			16'b100000000 : data = 16'b10111011;
			16'b100011010 : data = 16'b11000000;
			16'b100110011 : data = 16'b11000101;
			16'b101001101 : data = 16'b11001001;
			16'b101100110 : data = 16'b11001101;
			16'b110000000 : data = 16'b11010001;
			16'b110011010 : data = 16'b11010101;
			16'b110110011 : data = 16'b11011000;
			16'b111001101 : data = 16'b11011100;
			16'b111100110 : data = 16'b11011111;
			16'b1000000000 : data = 16'b11100001;
			16'b1000011010 : data = 16'b11100100;
			16'b1000110011 : data = 16'b11100110;
			16'b1001001101 : data = 16'b11101001;
			16'b1001100110 : data = 16'b11101011;
			16'b1010000000 : data = 16'b11101101;
			16'b1010011010 : data = 16'b11101110;
			16'b1010110011 : data = 16'b11110000;
			16'b1011001101 : data = 16'b11110001;
			16'b1011100110 : data = 16'b11110011;
			16'b1100000000 : data = 16'b11110100;
			16'b1100011010 : data = 16'b11110101;
			16'b1100110011 : data = 16'b11110110;
			16'b1101001101 : data = 16'b11110111;
			16'b1101100110 : data = 16'b11111000;
			16'b1110000000 : data = 16'b11111000;
			16'b1110011010 : data = 16'b11111001;
			16'b1110110011 : data = 16'b11111010;
			16'b1111001101 : data = 16'b11111010;
			16'b1111100110 : data = 16'b11111011;
			16'b10000000000 : data = 16'b11111011;
			16'b10000011010 : data = 16'b11111100;
			16'b10000110011 : data = 16'b11111100;
			16'b10001001101 : data = 16'b11111101;
			16'b10001100110 : data = 16'b11111101;
			16'b10010000000 : data = 16'b11111101;
			16'b10010011010 : data = 16'b11111101;
			16'b10010110011 : data = 16'b11111110;
			16'b10011001101 : data = 16'b11111110;
			16'b10011100110 : data = 16'b11111110;
			16'b10100000000 : data = 16'b11111110;
			16'b10100011010 : data = 16'b11111110;
			16'b10100110011 : data = 16'b11111111;
			16'b10101001101 : data = 16'b11111111;
			16'b10101100110 : data = 16'b11111111;
			16'b10110000000 : data = 16'b11111111;
			16'b10110011010 : data = 16'b11111111;
			16'b10110110011 : data = 16'b11111111;
			16'b10111001101 : data = 16'b11111111;
			16'b10111100110 : data = 16'b11111111;
			16'b11000000000 : data = 16'b11111111;
		endcase	
	end
	
endmodule
