module rom(addr,data);
	input [5:0] addr;
	output reg [15:0] data;
	
	//Look-up Table of Sigmoid (X >=0)
	always @ (addr) begin
		case(addr)
			6'b0 : data = 16'b10000000;
			6'b1 : data = 16'b10001000;
			6'b10 : data = 16'b10010000;
			6'b11 : data = 16'b10011000;
			6'b100 : data = 16'b10011111;
			6'b101 : data = 16'b10100111;
			6'b110 : data = 16'b10101110;
			6'b111 : data = 16'b10110101;
			6'b1000 : data = 16'b10111011;
			6'b1001 : data = 16'b11000001;
			6'b1010 : data = 16'b11000111;
			6'b1011 : data = 16'b11001100;
			6'b1100 : data = 16'b11010001;
			6'b1101 : data = 16'b11010110;
			6'b1110 : data = 16'b11011010;
			6'b1111 : data = 16'b11011110;
			6'b10000 : data = 16'b11100001;
			6'b10001 : data = 16'b11100101;
			6'b10010 : data = 16'b11101000;
			6'b10011 : data = 16'b11101010;
			6'b10100 : data = 16'b11101101;
			6'b10101 : data = 16'b11101111;
			6'b10110 : data = 16'b11110001;
			6'b10111 : data = 16'b11110010;
			6'b11000 : data = 16'b11110100;
			6'b11001 : data = 16'b11110101;
			6'b11010 : data = 16'b11110110;
			6'b11011 : data = 16'b11111000;
			6'b11100 : data = 16'b11111000;
			6'b11101 : data = 16'b11111001;
			6'b11110 : data = 16'b11111010;
			6'b11111 : data = 16'b11111011;
			6'b100000 : data = 16'b11111011;
			6'b100001 : data = 16'b11111100;
			6'b100010 : data = 16'b11111100;
			6'b100011 : data = 16'b11111101;
			6'b100100 : data = 16'b11111101;
			6'b100101 : data = 16'b11111110;
			6'b100110 : data = 16'b11111110;
			6'b100111 : data = 16'b11111110;
			6'b101000 : data = 16'b11111110;
			6'b101001 : data = 16'b11111110;
			6'b101010 : data = 16'b11111111;
			6'b101011 : data = 16'b11111111;
			6'b101100 : data = 16'b11111111;
			6'b101101 : data = 16'b11111111;
			6'b101110 : data = 16'b11111111;
			6'b101111 : data = 16'b11111111;
			6'b110000 : data = 16'b11111111;
		endcase	
	end
	
endmodule
