
module Top ( clk, reset, Done );
  input clk, reset;
  output Done;
  wire   N3637, n24401, n24402, n36946, n36947, n36948, n36949, n36950, n36951,
         n36952, n36953, n36954, n36955, n36956, n36957, n36958, n36959,
         n36960, n36961, n36962, n36963, n36964, n36965, n36966, n36967,
         n36968, n36969, n36970, n36984, n36985, n36986, n36987, n36988,
         n36989, n36990, n36991, n36992, n36993, n36994, n36995, n36996,
         n36997, n36998, n36999, n37000, n37001, n37002, n37003, n37004,
         n37005, n37006, n37007, n37008, n37009, n37010, n37011, n37012,
         n37013, n37014, n37015, n37016, n37017, n37018, n37019, n37020,
         n37021, n37022, n37023, n37024, n37025, n37026, n37027, n37028,
         n37029, n37030, n37031, n37032, n37033, n37034, n37035, n37036,
         n37037, n37038, n37039, n37040, n37041, n37042, n37043, n37044,
         n37045, n37046, n37047, n37048, n37049, n37050, n37051, n37052,
         n37053, n37054, n37055, n37056, n37057, n37058, n37059, n37060,
         n37061, n37062, n37063, n37064, n37065, n37066, n37067, n37068,
         n37069, n37070, n37071, n37072, n37073, n37074, n37075, n37076,
         n37077, n37078, n37079, n37080, n37081, n37082, n37083, n37084,
         n37085, n37086, n37087, n37088, n37089, n37090, n37091, n37092,
         n37093, n37094, n37095, n37096, n37097, n37098, n37099, n37100,
         n37101, n37102, n37103, n37104, n37105, n37106, n37107, n37108,
         n37109, n37110, n37111, n37112, n37113, n37114, n37115, n37116,
         n37117, n37118, n37119, n37120, n37121, n37122, n37123, n37124,
         n37125, n37126, n37127, n37128, n37129, n37130, n37131, n37132,
         n37133, n37134, n37135, n37136, n37137, n37138, n37139, n37140,
         n37141, n37142, n37143, n37144, n37145, n37146, n37147, n37148,
         n37149, n37150, n37151;
  wire   [3:0] inoutAddrQ;
  wire   [1:0] midAddrQ;
  wire   [11:0] wAddrQ;
  wire   [1:0] currentState;
  wire   [5:0] wrCounterQ;

  dp_1 \currentState_reg[0]  ( .ip(n36969), .ck(clk), .q(currentState[0]) );
  dp_1 \currentState_reg[1]  ( .ip(n36970), .ck(clk), .q(currentState[1]) );
  dp_1 \wAddrQ_reg[11]  ( .ip(n36956), .ck(clk), .q(wAddrQ[11]) );
  dp_1 roundQ_reg ( .ip(n36968), .ck(clk), .q(N3637) );
  dp_1 \wAddrQ_reg[0]  ( .ip(n36967), .ck(clk), .q(wAddrQ[0]) );
  dp_1 \wAddrQ_reg[1]  ( .ip(n36966), .ck(clk), .q(wAddrQ[1]) );
  dp_1 \wAddrQ_reg[2]  ( .ip(n36965), .ck(clk), .q(wAddrQ[2]) );
  dp_1 \wAddrQ_reg[3]  ( .ip(n36964), .ck(clk), .q(wAddrQ[3]) );
  dp_1 \wAddrQ_reg[4]  ( .ip(n36963), .ck(clk), .q(wAddrQ[4]) );
  dp_1 \wAddrQ_reg[5]  ( .ip(n36962), .ck(clk), .q(wAddrQ[5]) );
  dp_1 \wAddrQ_reg[6]  ( .ip(n36961), .ck(clk), .q(wAddrQ[6]) );
  dp_1 \wAddrQ_reg[7]  ( .ip(n36960), .ck(clk), .q(wAddrQ[7]) );
  dp_1 \wAddrQ_reg[8]  ( .ip(n36959), .ck(clk), .q(wAddrQ[8]) );
  dp_1 \wAddrQ_reg[9]  ( .ip(n36958), .ck(clk), .q(wAddrQ[9]) );
  dp_1 \wAddrQ_reg[10]  ( .ip(n36957), .ck(clk), .q(wAddrQ[10]) );
  dp_1 \wrCounterQ_reg[0]  ( .ip(n36955), .ck(clk), .q(wrCounterQ[0]) );
  dp_1 \wrCounterQ_reg[1]  ( .ip(n36954), .ck(clk), .q(wrCounterQ[1]) );
  dp_1 \wrCounterQ_reg[2]  ( .ip(n36953), .ck(clk), .q(wrCounterQ[2]) );
  dp_1 \wrCounterQ_reg[3]  ( .ip(n36952), .ck(clk), .q(wrCounterQ[3]) );
  dp_1 \wrCounterQ_reg[4]  ( .ip(n36951), .ck(clk), .q(wrCounterQ[4]) );
  dp_1 \wrCounterQ_reg[5]  ( .ip(n36950), .ck(clk), .q(wrCounterQ[5]) );
  dp_1 \midAddrQ_reg[1]  ( .ip(n24401), .ck(clk), .q(midAddrQ[1]) );
  dp_1 \midAddrQ_reg[0]  ( .ip(n24402), .ck(clk), .q(midAddrQ[0]) );
  dp_1 \inoutAddrQ_reg[0]  ( .ip(n36949), .ck(clk), .q(inoutAddrQ[0]) );
  dp_1 \inoutAddrQ_reg[3]  ( .ip(n36946), .ck(clk), .q(inoutAddrQ[3]) );
  dp_1 \inoutAddrQ_reg[1]  ( .ip(n36948), .ck(clk), .q(inoutAddrQ[1]) );
  dp_1 \inoutAddrQ_reg[2]  ( .ip(n36947), .ck(clk), .q(inoutAddrQ[2]) );
  inv_1 U38062 ( .ip(wrCounterQ[4]), .op(n37092) );
  inv_1 U38063 ( .ip(reset), .op(n37012) );
  inv_1 U38064 ( .ip(currentState[1]), .op(n37042) );
  nor2_1 U38065 ( .ip1(currentState[0]), .ip2(n37042), .op(n37131) );
  inv_1 U38066 ( .ip(n37131), .op(n37008) );
  nand2_1 U38067 ( .ip1(n37012), .ip2(n37008), .op(n37086) );
  inv_1 U38068 ( .ip(n37086), .op(n36997) );
  inv_1 U38069 ( .ip(N3637), .op(n37132) );
  nor4_1 U38070 ( .ip1(wAddrQ[4]), .ip2(wAddrQ[1]), .ip3(wAddrQ[2]), .ip4(
        wAddrQ[0]), .op(n36985) );
  inv_1 U38071 ( .ip(wAddrQ[6]), .op(n36984) );
  nand4_1 U38072 ( .ip1(wAddrQ[5]), .ip2(wAddrQ[3]), .ip3(n36985), .ip4(n36984), .op(n37010) );
  nor2_1 U38073 ( .ip1(wAddrQ[8]), .ip2(wAddrQ[7]), .op(n36989) );
  inv_1 U38074 ( .ip(wAddrQ[10]), .op(n37017) );
  nand4_1 U38075 ( .ip1(n36989), .ip2(wAddrQ[11]), .ip3(wAddrQ[9]), .ip4(
        n37017), .op(n37009) );
  nor2_1 U38076 ( .ip1(n37010), .ip2(n37009), .op(n36986) );
  nor2_1 U38077 ( .ip1(n36986), .ip2(n37008), .op(n37140) );
  nand3_1 U38078 ( .ip1(n37132), .ip2(n37140), .ip3(n37012), .op(n36991) );
  nand2_1 U38079 ( .ip1(N3637), .ip2(n37131), .op(n37011) );
  inv_1 U38080 ( .ip(n37011), .op(n37098) );
  inv_1 U38081 ( .ip(n37010), .op(n36990) );
  nor2_1 U38082 ( .ip1(wAddrQ[10]), .ip2(wAddrQ[9]), .op(n36988) );
  inv_1 U38083 ( .ip(wAddrQ[11]), .op(n36987) );
  nand4_1 U38084 ( .ip1(n36990), .ip2(n36989), .ip3(n36988), .ip4(n36987), 
        .op(n37041) );
  nand3_1 U38085 ( .ip1(n37098), .ip2(n37041), .ip3(n37012), .op(n37104) );
  nand2_1 U38086 ( .ip1(n36991), .ip2(n37104), .op(n37094) );
  nor2_1 U38087 ( .ip1(n36997), .ip2(n37094), .op(n36998) );
  nand3_1 U38088 ( .ip1(wrCounterQ[1]), .ip2(wrCounterQ[2]), .ip3(
        wrCounterQ[0]), .op(n37089) );
  inv_1 U38089 ( .ip(wrCounterQ[3]), .op(n37088) );
  nor2_1 U38090 ( .ip1(n37089), .ip2(n37088), .op(n37101) );
  and3_1 U38091 ( .ip1(n37086), .ip2(wrCounterQ[4]), .ip3(n37101), .op(n36992)
         );
  nor2_1 U38092 ( .ip1(n36998), .ip2(n36992), .op(n37095) );
  inv_1 U38093 ( .ip(n37095), .op(n36993) );
  or2_1 U38094 ( .ip1(n37092), .ip2(n36993), .op(n36996) );
  nand2_1 U38095 ( .ip1(n37101), .ip2(n37094), .op(n36994) );
  or2_1 U38096 ( .ip1(n36994), .ip2(n36993), .op(n36995) );
  nand2_1 U38097 ( .ip1(n36996), .ip2(n36995), .op(n36951) );
  inv_1 U38098 ( .ip(wrCounterQ[1]), .op(n37083) );
  or2_1 U38099 ( .ip1(wrCounterQ[1]), .ip2(n36998), .op(n37000) );
  inv_1 U38100 ( .ip(wrCounterQ[0]), .op(n37005) );
  nor2_1 U38101 ( .ip1(n36997), .ip2(n37005), .op(n37004) );
  or2_1 U38102 ( .ip1(n37004), .ip2(n36998), .op(n36999) );
  nand2_1 U38103 ( .ip1(n37000), .ip2(n36999), .op(n37084) );
  inv_1 U38104 ( .ip(n37084), .op(n37001) );
  or2_1 U38105 ( .ip1(n37083), .ip2(n37001), .op(n37003) );
  nand2_1 U38106 ( .ip1(wrCounterQ[0]), .ip2(n37094), .op(n37082) );
  or2_1 U38107 ( .ip1(n37082), .ip2(n37001), .op(n37002) );
  nand2_1 U38108 ( .ip1(n37003), .ip2(n37002), .op(n36954) );
  inv_1 U38109 ( .ip(n37094), .op(n37087) );
  or2_1 U38110 ( .ip1(n37087), .ip2(n37004), .op(n37007) );
  or2_1 U38111 ( .ip1(n37005), .ip2(n37004), .op(n37006) );
  nand2_1 U38112 ( .ip1(n37007), .ip2(n37006), .op(n36955) );
  nand2_1 U38113 ( .ip1(currentState[0]), .ip2(n37042), .op(n37144) );
  nor2_1 U38114 ( .ip1(reset), .ip2(n37144), .op(n37105) );
  or3_1 U38115 ( .ip1(n37010), .ip2(n37009), .ip3(n37008), .op(n37034) );
  nand4_1 U38116 ( .ip1(n37144), .ip2(n37012), .ip3(n37011), .ip4(n37034), 
        .op(n37013) );
  nand2_1 U38117 ( .ip1(n37104), .ip2(n37013), .op(n37072) );
  or2_1 U38118 ( .ip1(n37105), .ip2(n37072), .op(n37057) );
  inv_1 U38119 ( .ip(wAddrQ[4]), .op(n37030) );
  nand3_1 U38120 ( .ip1(wAddrQ[1]), .ip2(wAddrQ[2]), .ip3(wAddrQ[0]), .op(
        n37024) );
  inv_1 U38121 ( .ip(n37024), .op(n37014) );
  nand2_1 U38122 ( .ip1(wAddrQ[3]), .ip2(n37014), .op(n37055) );
  nor2_1 U38123 ( .ip1(n37030), .ip2(n37055), .op(n37028) );
  nand3_1 U38124 ( .ip1(wAddrQ[6]), .ip2(wAddrQ[5]), .ip3(n37028), .op(n37018)
         );
  or2_1 U38125 ( .ip1(n37018), .ip2(n37072), .op(n37015) );
  nand2_1 U38126 ( .ip1(n37057), .ip2(n37015), .op(n37067) );
  nand4_1 U38127 ( .ip1(wAddrQ[8]), .ip2(wAddrQ[7]), .ip3(wAddrQ[10]), .ip4(
        wAddrQ[9]), .op(n37078) );
  nand2_1 U38128 ( .ip1(n37105), .ip2(n37078), .op(n37016) );
  nand2_1 U38129 ( .ip1(n37067), .ip2(n37016), .op(n37080) );
  inv_1 U38130 ( .ip(n37080), .op(n37019) );
  or2_1 U38131 ( .ip1(n37017), .ip2(n37019), .op(n37022) );
  inv_1 U38132 ( .ip(wAddrQ[8]), .op(n37069) );
  inv_1 U38133 ( .ip(wAddrQ[7]), .op(n37068) );
  nor3_1 U38134 ( .ip1(n37069), .ip2(n37068), .ip3(n37018), .op(n37073) );
  nand3_1 U38135 ( .ip1(wAddrQ[9]), .ip2(n37105), .ip3(n37073), .op(n37020) );
  or2_1 U38136 ( .ip1(n37020), .ip2(n37019), .op(n37021) );
  nand2_1 U38137 ( .ip1(n37022), .ip2(n37021), .op(n36957) );
  nand2_1 U38138 ( .ip1(n37105), .ip2(n37068), .op(n37023) );
  nand2_1 U38139 ( .ip1(n37067), .ip2(n37023), .op(n37071) );
  inv_1 U38140 ( .ip(n37071), .op(n37025) );
  or2_1 U38141 ( .ip1(n37068), .ip2(n37025), .op(n37027) );
  inv_1 U38142 ( .ip(n37105), .op(n37049) );
  nor2_1 U38143 ( .ip1(n37049), .ip2(n37024), .op(n37058) );
  nand2_1 U38144 ( .ip1(wAddrQ[3]), .ip2(n37058), .op(n37031) );
  nor2_1 U38145 ( .ip1(n37030), .ip2(n37031), .op(n37063) );
  nand3_1 U38146 ( .ip1(wAddrQ[6]), .ip2(wAddrQ[5]), .ip3(n37063), .op(n37079)
         );
  or2_1 U38147 ( .ip1(n37079), .ip2(n37025), .op(n37026) );
  nand2_1 U38148 ( .ip1(n37027), .ip2(n37026), .op(n36960) );
  nor2_1 U38149 ( .ip1(n37028), .ip2(n37049), .op(n37029) );
  nor2_1 U38150 ( .ip1(n37029), .ip2(n37072), .op(n37061) );
  or2_1 U38151 ( .ip1(n37030), .ip2(n37061), .op(n37033) );
  or2_1 U38152 ( .ip1(n37031), .ip2(n37061), .op(n37032) );
  nand2_1 U38153 ( .ip1(n37033), .ip2(n37032), .op(n36963) );
  or2_1 U38154 ( .ip1(n37132), .ip2(reset), .op(n37036) );
  or2_1 U38155 ( .ip1(n37034), .ip2(reset), .op(n37035) );
  nand2_1 U38156 ( .ip1(n37036), .ip2(n37035), .op(n36968) );
  and2_1 U38157 ( .ip1(currentState[0]), .ip2(currentState[1]), .op(Done) );
  nand2_1 U38158 ( .ip1(midAddrQ[1]), .ip2(midAddrQ[0]), .op(n37148) );
  or3_1 U38159 ( .ip1(n37132), .ip2(n37148), .ip3(n37144), .op(n37040) );
  inv_1 U38160 ( .ip(inoutAddrQ[0]), .op(n37111) );
  inv_1 U38161 ( .ip(inoutAddrQ[1]), .op(n37037) );
  nand4_1 U38162 ( .ip1(n37111), .ip2(n37037), .ip3(inoutAddrQ[3]), .ip4(
        inoutAddrQ[2]), .op(n37107) );
  inv_1 U38163 ( .ip(n37107), .op(n37038) );
  nor2_1 U38164 ( .ip1(N3637), .ip2(n37144), .op(n37099) );
  nand2_1 U38165 ( .ip1(n37038), .ip2(n37099), .op(n37039) );
  nand2_1 U38166 ( .ip1(n37040), .ip2(n37039), .op(n37045) );
  nor3_1 U38167 ( .ip1(n37132), .ip2(n37042), .ip3(n37041), .op(n37043) );
  nor3_1 U38168 ( .ip1(Done), .ip2(n37045), .ip3(n37043), .op(n37044) );
  nor2_1 U38169 ( .ip1(reset), .ip2(n37044), .op(n36970) );
  nor2_1 U38170 ( .ip1(reset), .ip2(n37045), .op(n36969) );
  mux2_1 U38171 ( .ip1(n37105), .ip2(n37072), .s(wAddrQ[0]), .op(n36967) );
  nand2_1 U38172 ( .ip1(wAddrQ[1]), .ip2(n37072), .op(n37048) );
  or2_1 U38173 ( .ip1(wAddrQ[1]), .ip2(wAddrQ[0]), .op(n37046) );
  nand2_1 U38174 ( .ip1(wAddrQ[1]), .ip2(wAddrQ[0]), .op(n37050) );
  nand3_1 U38175 ( .ip1(n37105), .ip2(n37046), .ip3(n37050), .op(n37047) );
  nand2_1 U38176 ( .ip1(n37048), .ip2(n37047), .op(n36966) );
  nor2_1 U38177 ( .ip1(n37050), .ip2(n37049), .op(n37054) );
  inv_1 U38178 ( .ip(n37072), .op(n37052) );
  nand2_1 U38179 ( .ip1(n37050), .ip2(n37105), .op(n37051) );
  nand2_1 U38180 ( .ip1(n37052), .ip2(n37051), .op(n37053) );
  mux2_1 U38181 ( .ip1(n37054), .ip2(n37053), .s(wAddrQ[2]), .op(n36965) );
  or2_1 U38182 ( .ip1(n37055), .ip2(n37072), .op(n37056) );
  nand2_1 U38183 ( .ip1(n37057), .ip2(n37056), .op(n37060) );
  nor2_1 U38184 ( .ip1(wAddrQ[3]), .ip2(n37058), .op(n37059) );
  nor2_1 U38185 ( .ip1(n37060), .ip2(n37059), .op(n36964) );
  inv_1 U38186 ( .ip(n37061), .op(n37062) );
  mux2_1 U38187 ( .ip1(n37063), .ip2(n37062), .s(wAddrQ[5]), .op(n36962) );
  or2_1 U38188 ( .ip1(wAddrQ[5]), .ip2(wAddrQ[6]), .op(n37065) );
  or2_1 U38189 ( .ip1(n37063), .ip2(wAddrQ[6]), .op(n37064) );
  nand2_1 U38190 ( .ip1(n37065), .ip2(n37064), .op(n37066) );
  nor2_1 U38191 ( .ip1(n37067), .ip2(n37066), .op(n36961) );
  nor2_1 U38192 ( .ip1(n37068), .ip2(n37079), .op(n37070) );
  mux2_1 U38193 ( .ip1(n37071), .ip2(n37070), .s(n37069), .op(n36959) );
  nand2_1 U38194 ( .ip1(wAddrQ[9]), .ip2(n37072), .op(n37077) );
  inv_1 U38195 ( .ip(wAddrQ[9]), .op(n37074) );
  mux2_1 U38196 ( .ip1(wAddrQ[9]), .ip2(n37074), .s(n37073), .op(n37075) );
  nand2_1 U38197 ( .ip1(n37105), .ip2(n37075), .op(n37076) );
  nand2_1 U38198 ( .ip1(n37077), .ip2(n37076), .op(n36958) );
  nor2_1 U38199 ( .ip1(n37079), .ip2(n37078), .op(n37081) );
  mux2_1 U38200 ( .ip1(n37081), .ip2(n37080), .s(wAddrQ[11]), .op(n36956) );
  nor2_1 U38201 ( .ip1(n37083), .ip2(n37082), .op(n37085) );
  mux2_1 U38202 ( .ip1(n37085), .ip2(n37084), .s(wrCounterQ[2]), .op(n36953)
         );
  nor2_1 U38203 ( .ip1(n37088), .ip2(n37086), .op(n37091) );
  not_ab_or_c_or_d U38204 ( .ip1(n37089), .ip2(n37088), .ip3(n37087), .ip4(
        n37101), .op(n37090) );
  or2_1 U38205 ( .ip1(n37091), .ip2(n37090), .op(n36952) );
  nor2_1 U38206 ( .ip1(wrCounterQ[5]), .ip2(n37092), .op(n37093) );
  nand3_1 U38207 ( .ip1(n37094), .ip2(n37093), .ip3(n37101), .op(n37097) );
  nand2_1 U38208 ( .ip1(wrCounterQ[5]), .ip2(n37095), .op(n37096) );
  nand2_1 U38209 ( .ip1(n37097), .ip2(n37096), .op(n36950) );
  inv_1 U38210 ( .ip(n37104), .op(n37100) );
  nor3_1 U38211 ( .ip1(n37099), .ip2(reset), .ip3(n37098), .op(n37110) );
  or2_1 U38212 ( .ip1(n37100), .ip2(n37110), .op(n37103) );
  nand3_1 U38213 ( .ip1(n37101), .ip2(wrCounterQ[4]), .ip3(wrCounterQ[5]), 
        .op(n37139) );
  or2_1 U38214 ( .ip1(n37139), .ip2(n37110), .op(n37102) );
  nand2_1 U38215 ( .ip1(n37103), .ip2(n37102), .op(n37113) );
  inv_1 U38216 ( .ip(n37113), .op(n37116) );
  nor2_1 U38217 ( .ip1(n37139), .ip2(n37104), .op(n37106) );
  or2_1 U38218 ( .ip1(n37105), .ip2(n37106), .op(n37109) );
  or2_1 U38219 ( .ip1(n37107), .ip2(n37106), .op(n37108) );
  nand2_1 U38220 ( .ip1(n37109), .ip2(n37108), .op(n37115) );
  nor2_1 U38221 ( .ip1(n37110), .ip2(n37115), .op(n37125) );
  mux2_1 U38222 ( .ip1(n37116), .ip2(n37125), .s(n37111), .op(n36949) );
  and2_1 U38223 ( .ip1(inoutAddrQ[0]), .ip2(n37125), .op(n37120) );
  nand2_1 U38224 ( .ip1(n37125), .ip2(n37111), .op(n37112) );
  nand2_1 U38225 ( .ip1(n37113), .ip2(n37112), .op(n37114) );
  mux2_1 U38226 ( .ip1(n37120), .ip2(n37114), .s(inoutAddrQ[1]), .op(n36948)
         );
  nand3_1 U38227 ( .ip1(inoutAddrQ[0]), .ip2(inoutAddrQ[1]), .ip3(
        inoutAddrQ[2]), .op(n37124) );
  or2_1 U38228 ( .ip1(n37124), .ip2(n37116), .op(n37119) );
  inv_1 U38229 ( .ip(n37115), .op(n37117) );
  or2_1 U38230 ( .ip1(n37117), .ip2(n37116), .op(n37118) );
  nand2_1 U38231 ( .ip1(n37119), .ip2(n37118), .op(n37128) );
  or2_1 U38232 ( .ip1(inoutAddrQ[1]), .ip2(inoutAddrQ[2]), .op(n37122) );
  or2_1 U38233 ( .ip1(n37120), .ip2(inoutAddrQ[2]), .op(n37121) );
  nand2_1 U38234 ( .ip1(n37122), .ip2(n37121), .op(n37123) );
  nor2_1 U38235 ( .ip1(n37128), .ip2(n37123), .op(n36947) );
  nor2_1 U38236 ( .ip1(inoutAddrQ[3]), .ip2(n37124), .op(n37126) );
  nand2_1 U38237 ( .ip1(n37126), .ip2(n37125), .op(n37130) );
  inv_1 U38238 ( .ip(inoutAddrQ[3]), .op(n37127) );
  or2_1 U38239 ( .ip1(n37128), .ip2(n37127), .op(n37129) );
  nand2_1 U38240 ( .ip1(n37130), .ip2(n37129), .op(n36946) );
  nor2_1 U38241 ( .ip1(n37132), .ip2(n37144), .op(n37135) );
  nand2_1 U38242 ( .ip1(n37132), .ip2(n37131), .op(n37133) );
  inv_1 U38243 ( .ip(n37133), .op(n37134) );
  nor2_1 U38244 ( .ip1(n37135), .ip2(n37134), .op(n37142) );
  or2_1 U38245 ( .ip1(n37140), .ip2(n37142), .op(n37137) );
  or2_1 U38246 ( .ip1(n37139), .ip2(n37142), .op(n37136) );
  nand2_1 U38247 ( .ip1(n37137), .ip2(n37136), .op(n37138) );
  nor2_1 U38248 ( .ip1(reset), .ip2(n37138), .op(n37149) );
  inv_1 U38249 ( .ip(n37139), .op(n37141) );
  nand2_1 U38250 ( .ip1(n37141), .ip2(n37140), .op(n37143) );
  not_ab_or_c_or_d U38251 ( .ip1(n37144), .ip2(n37143), .ip3(n37142), .ip4(
        reset), .op(n37147) );
  inv_1 U38252 ( .ip(midAddrQ[0]), .op(n37145) );
  mux2_1 U38253 ( .ip1(n37149), .ip2(n37147), .s(n37145), .op(n24402) );
  or2_1 U38254 ( .ip1(midAddrQ[1]), .ip2(midAddrQ[0]), .op(n37146) );
  nand3_1 U38255 ( .ip1(n37148), .ip2(n37147), .ip3(n37146), .op(n37151) );
  nand2_1 U38256 ( .ip1(midAddrQ[1]), .ip2(n37149), .op(n37150) );
  nand2_1 U38257 ( .ip1(n37151), .ip2(n37150), .op(n24401) );
endmodule

