module rom(addr,data)
	input [6:0] addr;
	output reg [15:0] data;
	
	//Look-up Table of Sigmoid
	always @ (addr) begin
		case(addr)
			16'b1111101000000000 : data = 16'b1;
			16'b1111101000011010 : data = 16'b1;
			16'b1111101000110010 : data = 16'b1;
			16'b1111101001001100 : data = 16'b1;
			16'b1111101001100110 : data = 16'b1;
			16'b1111101010000000 : data = 16'b1;
			16'b1111101010011010 : data = 16'b1;
			16'b1111101010110010 : data = 16'b1;
			16'b1111101011001100 : data = 16'b1;
			16'b1111101011100110 : data = 16'b10;
			16'b1111101100000000 : data = 16'b10;
			16'b1111101100011010 : data = 16'b10;
			16'b1111101100110010 : data = 16'b10;
			16'b1111101101001100 : data = 16'b10;
			16'b1111101101100110 : data = 16'b11;
			16'b1111101110000000 : data = 16'b11;
			16'b1111101110011010 : data = 16'b11;
			16'b1111101110110010 : data = 16'b11;
			16'b1111101111001100 : data = 16'b100;
			16'b1111101111100110 : data = 16'b100;
			16'b1111110000000000 : data = 16'b101;
			16'b1111110000011010 : data = 16'b101;
			16'b1111110000110010 : data = 16'b110;
			16'b1111110001001100 : data = 16'b110;
			16'b1111110001100110 : data = 16'b111;
			16'b1111110010000000 : data = 16'b1000;
			16'b1111110010011010 : data = 16'b1000;
			16'b1111110010110010 : data = 16'b1001;
			16'b1111110011001100 : data = 16'b1010;
			16'b1111110011100110 : data = 16'b1011;
			16'b1111110100000000 : data = 16'b1100;
			16'b1111110100011010 : data = 16'b1101;
			16'b1111110100110010 : data = 16'b1111;
			16'b1111110101001100 : data = 16'b10000;
			16'b1111110101100110 : data = 16'b10010;
			16'b1111110110000000 : data = 16'b10011;
			16'b1111110110011010 : data = 16'b10101;
			16'b1111110110110010 : data = 16'b10111;
			16'b1111110111001100 : data = 16'b11010;
			16'b1111110111100110 : data = 16'b11100;
			16'b1111111000000000 : data = 16'b11111;
			16'b1111111000011010 : data = 16'b100001;
			16'b1111111000110010 : data = 16'b100100;
			16'b1111111001001100 : data = 16'b101000;
			16'b1111111001100110 : data = 16'b101011;
			16'b1111111010000000 : data = 16'b101111;
			16'b1111111010011010 : data = 16'b110011;
			16'b1111111010110010 : data = 16'b110111;
			16'b1111111011001100 : data = 16'b111011;
			16'b1111111011100110 : data = 16'b1000000;
			16'b1111111100000000 : data = 16'b1000101;
			16'b1111111100011010 : data = 16'b1001010;
			16'b1111111100110010 : data = 16'b1001111;
			16'b1111111101001100 : data = 16'b1010101;
			16'b1111111101100110 : data = 16'b1011011;
			16'b1111111110000000 : data = 16'b1100001;
			16'b1111111110011010 : data = 16'b1100111;
			16'b1111111110110010 : data = 16'b1101101;
			16'b1111111111001100 : data = 16'b1110011;
			16'b1111111111100110 : data = 16'b1111010;
			16'b0 : data = 16'b10000000;
			16'b11010 : data = 16'b10000110;
			16'b110011 : data = 16'b10001101;
			16'b1001101 : data = 16'b10010011;
			16'b1100110 : data = 16'b10011001;
			16'b10000000 : data = 16'b10011111;
			16'b10011010 : data = 16'b10100101;
			16'b10110011 : data = 16'b10101011;
			16'b11001101 : data = 16'b10110001;
			16'b11100110 : data = 16'b10110110;
			16'b100000000 : data = 16'b10111011;
			16'b100011010 : data = 16'b11000000;
			16'b100110011 : data = 16'b11000101;
			16'b101001101 : data = 16'b11001001;
			16'b101100110 : data = 16'b11001101;
			16'b110000000 : data = 16'b11010001;
			16'b110011010 : data = 16'b11010101;
			16'b110110011 : data = 16'b11011000;
			16'b111001101 : data = 16'b11011100;
			16'b111100110 : data = 16'b11011111;
			16'b1000000000 : data = 16'b11100001;
			16'b1000011010 : data = 16'b11100100;
			16'b1000110011 : data = 16'b11100110;
			16'b1001001101 : data = 16'b11101001;
			16'b1001100110 : data = 16'b11101011;
			16'b1010000000 : data = 16'b11101101;
			16'b1010011010 : data = 16'b11101110;
			16'b1010110011 : data = 16'b11110000;
			16'b1011001101 : data = 16'b11110001;
			16'b1011100110 : data = 16'b11110011;
			16'b1100000000 : data = 16'b11110100;
			16'b1100011010 : data = 16'b11110101;
			16'b1100110011 : data = 16'b11110110;
			16'b1101001101 : data = 16'b11110111;
			16'b1101100110 : data = 16'b11111000;
			16'b1110000000 : data = 16'b11111000;
			16'b1110011010 : data = 16'b11111001;
			16'b1110110011 : data = 16'b11111010;
			16'b1111001101 : data = 16'b11111010;
			16'b1111100110 : data = 16'b11111011;
			16'b10000000000 : data = 16'b11111011;
			16'b10000011010 : data = 16'b11111100;
			16'b10000110011 : data = 16'b11111100;
			16'b10001001101 : data = 16'b11111101;
			16'b10001100110 : data = 16'b11111101;
			16'b10010000000 : data = 16'b11111101;
			16'b10010011010 : data = 16'b11111101;
			16'b10010110011 : data = 16'b11111110;
			16'b10011001101 : data = 16'b11111110;
			16'b10011100110 : data = 16'b11111110;
			16'b10100000000 : data = 16'b11111110;
			16'b10100011010 : data = 16'b11111110;
			16'b10100110011 : data = 16'b11111111;
			16'b10101001101 : data = 16'b11111111;
			16'b10101100110 : data = 16'b11111111;
			16'b10110000000 : data = 16'b11111111;
			16'b10110011010 : data = 16'b11111111;
			16'b10110110011 : data = 16'b11111111;
			16'b10111001101 : data = 16'b11111111;
			16'b10111100110 : data = 16'b11111111;
			16'b11000000000 : data = 16'b11111111;
		endcase	
	end
	
endmodule
